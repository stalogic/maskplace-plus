version https://git-lfs.github.com/spec/v1
oid sha256:9bda2ceb1151dc9cdf0f14a514658a91b561681783d232e1badad1fdfcdd92aa
size 15333
