version https://git-lfs.github.com/spec/v1
oid sha256:834a79295054cd4209178d1bade67c353863c47bb4b3c22ee38b862b7cec37f2
size 19485
