version https://git-lfs.github.com/spec/v1
oid sha256:2a5df0db471b7b824e9052fadbe11ee64ea1ecfc549a43df0e8941b90e607de4
size 326014
