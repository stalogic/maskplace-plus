version https://git-lfs.github.com/spec/v1
oid sha256:ae48ca01bc12b9f0c44717b7275ba8884f1760bf562f5a42e3ca39906ddc9e54
size 255850
